`ifndef SCOREBOARD_V
`define SCOREBOARD_V

module Scoreboard (
    input            clock,
    input            reset,

    // Issue stage asynchronous read interface
    input      [4:0] iss_ass_addr_a,      // requested register
    output           iss_ass_pending_a,   // register status
    output     [1:0] iss_ass_unit_a,      // register functional unit
    output     [4:0] iss_ass_row_a,       // register execution stage

    input      [4:0] iss_ass_addr_b,      // requested register
    output           iss_ass_pending_b,   // register status
    output     [1:0] iss_ass_unit_b,      // register functional unit
    output     [4:0] iss_ass_row_b,       // register execution stage

    // Decode stage asynchronous read interface
    input      [4:0] id_ass_addr_a,      // requested register
    output           id_ass_pending_a,   // register status
    output     [1:0] id_ass_unit_a,      // register functional unit
    output     [4:0] id_ass_row_a,       // register execution stage

    input      [4:0] id_ass_addr_b,      // requested register
    output           id_ass_pending_b,   // register status
    output     [1:0] id_ass_unit_b,      // register functional unit
    output     [4:0] id_ass_row_b,       // register execution stage

    // Issue stage synchronous write interface
    input      [4:0] writeaddr,     // register to become pending
    input      [1:0] registerunit,  // which functional unit it is going to
    // 2'b00: AluMisc
    // 2'b01: Mem
    // 2'b10: Mult
    input            enablewrite   // prevent incorrect write (e.g. during stalls)
);

    reg [7:0] rows[31:0];
    reg [5:0] i;

    // outputs requested register data
    assign iss_ass_pending_a = rows[iss_ass_addr_a][7];
    assign iss_ass_unit_a    = rows[iss_ass_addr_a][6:5];
    assign iss_ass_row_a     = rows[iss_ass_addr_a][4:0];

    assign iss_ass_pending_b = rows[iss_ass_addr_b][7];
    assign iss_ass_unit_b    = rows[iss_ass_addr_b][6:5];
    assign iss_ass_row_b     = rows[iss_ass_addr_b][4:0];

    assign id_ass_pending_a = rows[id_ass_addr_a][7];
    assign id_ass_unit_a    = rows[id_ass_addr_a][6:5];
    assign id_ass_row_a     = rows[id_ass_addr_a][4:0];

    assign id_ass_pending_b = rows[id_ass_addr_b][7];
    assign id_ass_unit_b    = rows[id_ass_addr_b][6:5];
    assign id_ass_row_b     = rows[id_ass_addr_b][4:0];

    always @(posedge clock or negedge reset) begin
        if(~reset) begin

            for (i=0; i<32; i=i+1) begin
                rows[i] <= 8'b0ZZ00000;
            end

        end else begin

            for (i=0; i<32; i=i+1) begin
                // updates the positions of the data
                rows[i][4:0] = rows[i][4:0] >> 1;
                if(rows[i][4:0] == 5'b00000) begin
                    // register is not pending anymore
                    rows[i][7:5] = 3'b0ZZ;
                end
            end

            // writes registers claimed on issue stage
            if(enablewrite) begin
                // the corresponding register becomes pending
                // and we write its functional unity
                rows[writeaddr][7] = 1'b1;
                rows[writeaddr][6:5] = registerunit;
                case (registerunit)
                    2'b00: rows[writeaddr][1] = 1'b1; // am
                    2'b01: rows[writeaddr][2] = 1'b1; // mem
                    2'b10: rows[writeaddr][4] = 1'b1; // mult
                    // The two below should hopefully never happen
                    2'b11: rows[writeaddr][4] = 1'b1;
                    default: rows[writeaddr][4] = 1'b1;
                endcase
            end

        end
    end

endmodule

`endif
