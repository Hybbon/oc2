`ifndef HAZARDDETECTOR_V
`define HAZARDDETECTOR_V

module HazardDetector (
    input [4:0] rega,
    input [4:0] regb,
    
    output stalled 
);



endmodule

`endif